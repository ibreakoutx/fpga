library verilog;
use verilog.vl_types.all;
entity hfifo_stim_test is
end hfifo_stim_test;
